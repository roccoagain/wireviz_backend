* RC Low-Pass Filter Netlist for ngspice

* Input source with AC amplitude = 1 V
Vin in 0 AC 1

* Low-pass filter: R in series, C to ground
R1 in out 1k
C1 out 0 1uF

.control
  * Perform an AC analysis from 10 Hz to 100 MHz in decade steps
  ac dec 100 10 100MEG
  
  * Write frequency response data to CSV
  wrdata rc_lpf_data.csv frequency vdb(out) vp(out)
.endc

.end
